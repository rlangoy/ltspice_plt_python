*OPA314 (PSpice format)


* OPA314 SIMULATION MODEL
********************************************

* GREEN-LIS MACROMODEL ARCHITECTURE

********************************************
**  THIS FILE WAS CREATED BY TINA      **
**    (C) 1996-2006 DESIGNSOFT, INC.   **
********************************************


* REV A BY MAREK LIS; AUGUST 29, 2011
*
*
* THIS MACROMODEL HAS BEEN OPTIMIZED TO MODEL THE AC, DC, NOISE, AND TRANSIENT RESPONSE PERFORMANCE WITHIN 
* THE DEVICE DATA SHEET SPECIFIED LIMITS. CORRECT OPERATION OF THIS MACROMODEL HAS BEEN VERIFIED ON DESIGNSOFT
* TINA VERSION 7.0.80.224 SF. FOR HELP WITH OTHER ANALOG SIMULATION SOFTWARE, PLEASE CONSULT THE SOFTWARE SUPPLIER.
*
*  
* COPYRIGHT 2011 BY TEXAS INSTRUMENTS CORPORATION

* BEGIN MODEL OPA314

*GREEN-LIS MACRO-MODEL SIMULATED FEATURES:

*OPEN LOOP GAIN AND PHASE VS FREQUENCY WITH RL AND CL EFFECTS
*INPUT COMMON MODE REJECTION WITH FREQUENCY
*POWER SUPPLY REJECTION WITH FREQUENCY
*INPUT IMPEDANCE VS FREQUENCY 
*OUTPUT IMPEDANCE VS OUTPUT CURRENT
*INPUT VOLTAGE NOISE VS FREQUENCY
*INPUT CURRENT NOISE VS FREQUENCY 
*OUTPUT VOLTAGE SWING VS OUTPUT CURRENT
*SHORT-CIRCUIT OUTPUT CURRENT
*QUIESCENT CURRENT VS SUPPLY VOLTAGE
*SETTLING TIME VS CAPACITIVE LOAD
*SLEW RATE
*SMALL SIGNAL OVERSHOOT VS CAPACITIVE LOAD
*LARGE SIGNAL RESPONSE
*OVERLOAD RECOVERY TIME
*INPUT BIAS CURRENT
*INPUT VOLTAGE OFFSET
*INPUT COMMON MODE RANGE
*OUTPUT CURRENT COMING THROUGH THE SUPPLY RAILS

* PIN ORDER: +IN, -IN, V+, V-, OUT
.SUBCKT OPA314  1 2 3 4 5
V7          48 10 0
VOS         26 39 -375.1U
V11         52 53 100M
V10         54 55 100M
V6          9 60 10
V5          61 9 10
V4          57 59 7.8
V1          58 56 7.8
V9          72 11 0
IS2         3 26 400F
IS1         3 4 150U
IS3         44 4 -200F
V3          76 9 20
V2          9 77 20
R3          27 28 1MEG 
L4          9 28 17M IC=0 
XU15        12 9 29 30 VC_RES_0
L1          31 9 1F IC=0 
R2          31 32 1 
GVCCS8      9 32 9 33  1
XR109       34 9 RNOISE_FREE_0
C3          34 9 12F 
GVCCS4      9 34 23 9  1U
C2          35 9 5F 
XR109_2     35 9 RNOISE_FREE_1
GVCCS3      9 35 34 9  1M
R4          36 20 10M 
C7          37 38 1P 
C8          38 9 5P
CINNCM      9 37 5P 
XIN11       39 37 FEMT_0
L2          40 9 1F 
XR109_3     23 9 RNOISE_FREE_0
XR109_4     41 9 RNOISE_FREE_0
XVN11       38 39 VNSE_0
XU14        42 9 43 44 VCVS_LIMIT_0
L3          45 9 3.16M 
R1          40 42 1 
GVCCS2      9 42 9 46  1
XU13        10 47 IDEAL_D_0
EVCVS5      48 9 4 9  1
C11         41 9 12F
XR109_5     22 9 RNOISE_FREE_1
GVCCS12     9 23 41 9  1U
XU5         12 9 3 13 VCVS_LIMIT_1
XU6         9 12 14 4 VCVS_LIMIT_2
C15         3 4 10P IC=0 
C22         9 19 1P 
R29         19 21 1 
C23         9 24 1P IC=0 
C9          49 9 10P IC=0 
R26         49 12 10 
C21         9 15 1P IC=0 
C20         9 16 1P IC=0 
C19         17 9 1P IC=0 
C17         18 9 1P IC=0 
C16         9 50 1P IC=0 
C12         51 9 1P IC=0 
R13         30 24 1 
R36         24 55 1M 
R35         24 53 1M 
SW12        56 52 17 9  S_VSWITCH_1
SW11        54 57 9 18  S_VSWITCH_2
R34         24 58 1K 
R33         24 59 1K 
SW10        61 21 19 9  S_VSWITCH_3
SW9         21 60 9 19  S_VSWITCH_4
R25         62 17 1 
R19         63 18 1 
R16         64 50 1 
R14         65 51 1 
R12         66 15 1 
R7          67 16 1 
R5          68 22 10M 
R6          69 21 10M 
R15         0 9 100MEG 
C13         22 9 5F 
GVCCS1      9 22 35 9  1M
GISINKING   4 9 70 9  1M
GISOURCING  3 9 71 9  1M
R23         70 9 10K 
SW7         12 70 49 9  S_VSWITCH_5
R21         9 71 10K 
SW8         12 71 49 9  S_VSWITCH_6
SW4         69 66 15 9  S_VSWITCH_7
SW3         67 69 9 16  S_VSWITCH_8
XU3         57 25 67 9 VCVS_LIMIT_3
XU1         56 25 66 9 VCVS_LIMIT_3
SW2         36 62 17 9  S_VSWITCH_9
SW1         63 36 9 18  S_VSWITCH_10
XU8         26 3 IDEAL_D_1
XU12        4 26 IDEAL_D_1
EVCVS6      72 9 3 9  1
R22         73 47 100 
EVCVS4      73 9 26 9  1
XU2         47 11 IDEAL_D_0
SW6         68 64 50 9  S_VSWITCH_11
SW5         65 68 9 51  S_VSWITCH_12
XU26        47 44 9 74 VCCS_LIMIT_0
XU4         74 9 9 21 VCCS_LIMIT_1
LPSR        75 9 1M IC=0 
XVCVSPSRR   32 9 43 37 VCVS_LIMIT_4
XU22        76 12 63 9 VCVS_LIMIT_5
XU21        77 12 62 9 VCVS_LIMIT_5
XU20        14 5 64 9 VCVS_LIMIT_5
XU19        13 5 65 9 VCVS_LIMIT_6
XU11        4 44 IDEAL_D_1
XU10        44 3 IDEAL_D_1
C10         20 9 5F 
C5          23 9 12F 
XR109_6     20 9 RNOISE_FREE_1
GVCCS15     9 20 22 9  1M
GVCCS10     9 41 27 9  1U
R20         1 38 100 
R18         2 37 100 
GVCCS6      9 27 25 9  1U
XR102       78 79 RNOISE_FREE_0
XR101       80 78 RNOISE_FREE_0
C6          78 0 1 IC=0 
XR105       25 9 RNOISE_FREE_0
XR104       21 9 RNOISE_FREE_2
XR103       9 74 RNOISE_FREE_0
EVCVS34     9 0 78 0  1
RPSR        75 33 1 
GVCCS11     9 33 3 4  25U
RCM         45 46 1 
EVCVS29     80 0 3 0  1
EVCVS28     79 0 4 0  1
GVCCS7      9 46 26 9  15U
VCCVS1_IN   29 5
HCCVS1      12 9 VCCVS1_IN   1K
GVCCS5      9 25 21 9  1U
CCC         21 9 16U 
EVCVS3      30 9 20 9  1
.MODEL S_VSWITCH_1 VSWITCH (RON=1 ROFF=10MEG VON=100M VOFF=-100M)
.MODEL S_VSWITCH_2 VSWITCH (RON=1 ROFF=10MEG VON=100M VOFF=-100M)
.MODEL S_VSWITCH_3 VSWITCH (RON=10M ROFF=100MEG VON=150 VOFF=130)
.MODEL S_VSWITCH_4 VSWITCH (RON=10M ROFF=100MEG VON=150 VOFF=130)
.MODEL S_VSWITCH_5 VSWITCH (RON=1M ROFF=10MEG VON=-10M VOFF=0)
.MODEL S_VSWITCH_6 VSWITCH (RON=1M ROFF=10MEG VON=10M VOFF=0)
.MODEL S_VSWITCH_7 VSWITCH (RON=1 ROFF=10MEG VON=1 VOFF=-1)
.MODEL S_VSWITCH_8 VSWITCH (RON=1 ROFF=10MEG VON=1 VOFF=-1)
.MODEL S_VSWITCH_9 VSWITCH (RON=1 ROFF=1G VON=10 VOFF=-10)
.MODEL S_VSWITCH_10 VSWITCH (RON=1 ROFF=1G VON=10 VOFF=-10)
.MODEL S_VSWITCH_11 VSWITCH (RON=1 ROFF=1G VON=10 VOFF=-10)
.MODEL S_VSWITCH_12 VSWITCH (RON=1 ROFF=1G VON=10 VOFF=-10)
.ENDS


*VOLTAGE CONTROLLED RESISTOR
.SUBCKT VC_RES_0  1      2      3    4
*              VC+    VC-   RES1 RES2
*ERES 3 40 VALUE = {600*(I(VSENSE) /(1+ABS(V(1,2)))*0.075)}
ERES 3 40 VALUE = {600*(I(VSENSE) / SQRT(((ABS(V(1,2))/0.075)+1)/1))}
VSENSE 40 4 DC 0
.ENDS VC_RES_0 


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_0  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=1E6
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_0 


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_1  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=1E3
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_1 


* BEGIN PROG NSE FEMTO AMP/RT-HZ 
.SUBCKT FEMT_0  1 2
* BEGIN SETUP OF NOISE GEN - FEMPTOAMPS/RT-HZ
* INPUT THREE VARIABLES
* SET UP INSE 1/F
* FA/RHZ AT 1/F FREQ
.PARAM NLFF=5
* FREQ FOR 1/F VAL
.PARAM FLWF=0.001
* SET UP INSE FB
* FA/RHZ FLATBAND
.PARAM NVRF=5
* END USER INPUT
* START CALC VALS
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
* END CALC VALS
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
C1 1 0 1E-15
C2 2 0 1E-15
C3 1 2 1E-15
.ENDS
* END PROG NSE FEMTO AMP/RT-HZ


* BEGIN PROG NSE NANO VOLT/RT-HZ
.SUBCKT VNSE_0  1 2
* BEGIN SETUP OF NOISE GEN - NANOVOLT/RT-HZ
* INPUT THREE VARIABLES
* SET UP VNSE 1/F
* NV/RHZ AT 1/F FREQ
.PARAM NLF=150
* FREQ FOR 1/F VAL
.PARAM FLW=1
* SET UP VNSE FB
* NV/RHZ FLATBAND
.PARAM NVR=13
* END USER INPUT
* START CALC VALS
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
* END CALC VALS
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
C1 1 0 1E-15
C2 2 0 1E-15
C3 1 2 1E-15
.ENDS
* END PROG NSE NANOV/RT-HZ


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_0  VC+ VC- VOUT+ VOUT-
*              
.PARAM GAIN = 1
.PARAM VPOS = 10M
.PARAM VNEG = -10M
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VNEG,VPOS)}
.ENDS VCVS_LIMIT_0 


*TG IDEAL DIODE
.SUBCKT IDEAL_D_0  A C
D1 A C DNOM
.MODEL DNOM D (TT=10P CJO=1E-18 IS=1E-15 RS=1E-3)
.ENDS IDEAL_D_0 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_1  VC+ VC- VOUT+ VOUT-
*              

E1 VOUT+ VOUT- TABLE {ABS(V(VC+,VC-))} = (0,0.029) (0.25,0.029) (19.9,0.6) 
.ENDS VCVS_LIMIT_1 



*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_2  VC+ VC- VOUT+ VOUT-
*              

E1 VOUT+ VOUT- TABLE {ABS(V(VC+,VC-))} = (0,0.029) (0.25,0.029) (19.9,0.6)
.ENDS VCVS_LIMIT_2 



*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_3  VC+ VC- VOUT+ VOUT-
*              
.PARAM GAIN = 100
.PARAM VPOS = 6000
.PARAM VNEG = -6000
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VNEG,VPOS)}
.ENDS VCVS_LIMIT_3 


*TG IDEAL DIODE
.SUBCKT IDEAL_D_1  A C
D1 A C DNOM 
.MODEL DNOM D (TT=10P CJO=1E-18 IS=1E-15 RS=1E-3)
.ENDS IDEAL_D_1 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCCS_LIMIT_0  VC+ VC- IOUT+ IOUT-
*              
.PARAM GAIN = 100U
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS VCCS_LIMIT_0 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCCS_LIMIT_1  VC+ VC- IOUT+ IOUT-
*              
.PARAM GAIN = 3.25
.PARAM IPOS = 24
.PARAM INEG = -24
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS VCCS_LIMIT_1 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_4  VC+ VC- VOUT+ VOUT-
*              
.PARAM GAIN = -1
.PARAM VPOS = 10M
.PARAM VNEG = -10M
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VNEG,VPOS)}
.ENDS VCVS_LIMIT_4 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_5  VC+ VC- VOUT+ VOUT-
*              
.PARAM GAIN = 100
.PARAM VPOS = 5000
.PARAM VNEG = -5000
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VNEG,VPOS)}
.ENDS VCVS_LIMIT_5 


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_6  VC+ VC- VOUT+ VOUT-
*             
.PARAM GAIN = 100
.PARAM VPOS = 5000
.PARAM VNEG = -5000
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VNEG,VPOS)}
.ENDS VCVS_LIMIT_6 


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_2  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=3.16E3
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_2 


.END


.END
